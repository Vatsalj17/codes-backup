module and_module (
    a,
    b,
    c
);
  input a, b;
  output c;
  // assign c = a & b;
  and (c, a, b); // and(output, inputs)
endmodule
